// sll32_case.v
`timescale 1ns/1ps
module sll32(
    input  wire [31:0] a,
    input  wire [4:0]  shamt,
    output reg  [31:0] y
);
    always @(*) begin
        case (shamt)
            5'd0:  y = a;
            5'd1:  y = {a[30:0],  1'b0};
            5'd2:  y = {a[29:0],  2'b0};
            5'd3:  y = {a[28:0],  3'b0};
            5'd4:  y = {a[27:0],  4'b0};
            5'd5:  y = {a[26:0],  5'b0};
            5'd6:  y = {a[25:0],  6'b0};
            5'd7:  y = {a[24:0],  7'b0};
            5'd8:  y = {a[23:0],  8'b0};
            5'd9:  y = {a[22:0],  9'b0};
            5'd10: y = {a[21:0], 10'b0};
            5'd11: y = {a[20:0], 11'b0};
            5'd12: y = {a[19:0], 12'b0};
            5'd13: y = {a[18:0], 13'b0};
            5'd14: y = {a[17:0], 14'b0};
            5'd15: y = {a[16:0], 15'b0};
            5'd16: y = {a[15:0], 16'b0};
            5'd17: y = {a[14:0], 17'b0};
            5'd18: y = {a[13:0], 18'b0};
            5'd19: y = {a[12:0], 19'b0};
            5'd20: y = {a[11:0], 20'b0};
            5'd21: y = {a[10:0], 21'b0};
            5'd22: y = {a[9:0],  22'b0};
            5'd23: y = {a[8:0],  23'b0};
            5'd24: y = {a[7:0],  24'b0};
            5'd25: y = {a[6:0],  25'b0};
            5'd26: y = {a[5:0],  26'b0};
            5'd27: y = {a[4:0],  27'b0};
            5'd28: y = {a[3:0],  28'b0};
            5'd29: y = {a[2:0],  29'b0};
            5'd30: y = {a[1:0],  30'b0};
            5'd31: y = {a[0],    31'b0};
            default: y = 32'b0;
        endcase
    end
endmodule


// srl32_case.v
`timescale 1ns/1ps
module srl32 (
    input  wire [31:0] a,
    input  wire [4:0]  shamt,
    output reg  [31:0] y
);
    always @(*) begin
        case (shamt)
            5'd0:  y = a;
            5'd1:  y = {1'b0,        a[31:1]};
            5'd2:  y = {2'b0,        a[31:2]};
            5'd3:  y = {3'b0,        a[31:3]};
            5'd4:  y = {4'b0,        a[31:4]};
            5'd5:  y = {5'b0,        a[31:5]};
            5'd6:  y = {6'b0,        a[31:6]};
            5'd7:  y = {7'b0,        a[31:7]};
            5'd8:  y = {8'b0,        a[31:8]};
            5'd9:  y = {9'b0,        a[31:9]};
            5'd10: y = {10'b0,       a[31:10]};
            5'd11: y = {11'b0,       a[31:11]};
            5'd12: y = {12'b0,       a[31:12]};
            5'd13: y = {13'b0,       a[31:13]};
            5'd14: y = {14'b0,       a[31:14]};
            5'd15: y = {15'b0,       a[31:15]};
            5'd16: y = {16'b0,       a[31:16]};
            5'd17: y = {17'b0,       a[31:17]};
            5'd18: y = {18'b0,       a[31:18]};
            5'd19: y = {19'b0,       a[31:19]};
            5'd20: y = {20'b0,       a[31:20]};
            5'd21: y = {21'b0,       a[31:21]};
            5'd22: y = {22'b0,       a[31:22]};
            5'd23: y = {23'b0,       a[31:23]};
            5'd24: y = {24'b0,       a[31:24]};
            5'd25: y = {25'b0,       a[31:25]};
            5'd26: y = {26'b0,       a[31:26]};
            5'd27: y = {27'b0,       a[31:27]};
            5'd28: y = {28'b0,       a[31:28]};
            5'd29: y = {29'b0,       a[31:29]};
            5'd30: y = {30'b0,       a[31:30]};
            5'd31: y = {31'b0,       a[31]};
            default: y = 32'b0;
        endcase
    end
endmodule

// sra32_case.v
`timescale 1ns/1ps
module sra32 (
    input  wire [31:0] a,
    input  wire [4:0]  shamt,
    output reg  [31:0] y
);
    wire sign = a[31];
    always @(*) begin
        case (shamt)
            5'd0:  y = a;
            5'd1:  y = { {1{sign}},  a[31:1] };
            5'd2:  y = { {2{sign}},  a[31:2] };
            5'd3:  y = { {3{sign}},  a[31:3] };
            5'd4:  y = { {4{sign}},  a[31:4] };
            5'd5:  y = { {5{sign}},  a[31:5] };
            5'd6:  y = { {6{sign}},  a[31:6] };
            5'd7:  y = { {7{sign}},  a[31:7] };
            5'd8:  y = { {8{sign}},  a[31:8] };
            5'd9:  y = { {9{sign}},  a[31:9] };
            5'd10: y = { {10{sign}}, a[31:10]};
            5'd11: y = { {11{sign}}, a[31:11]};
            5'd12: y = { {12{sign}}, a[31:12]};
            5'd13: y = { {13{sign}}, a[31:13]};
            5'd14: y = { {14{sign}}, a[31:14]};
            5'd15: y = { {15{sign}}, a[31:15]};
            5'd16: y = { {16{sign}}, a[31:16]};
            5'd17: y = { {17{sign}}, a[31:17]};
            5'd18: y = { {18{sign}}, a[31:18]};
            5'd19: y = { {19{sign}}, a[31:19]};
            5'd20: y = { {20{sign}}, a[31:20]};
            5'd21: y = { {21{sign}}, a[31:21]};
            5'd22: y = { {22{sign}}, a[31:22]};
            5'd23: y = { {23{sign}}, a[31:23]};
            5'd24: y = { {24{sign}}, a[31:24]};
            5'd25: y = { {25{sign}}, a[31:25]};
            5'd26: y = { {26{sign}}, a[31:26]};
            5'd27: y = { {27{sign}}, a[31:27]};
            5'd28: y = { {28{sign}}, a[31:28]};
            5'd29: y = { {29{sign}}, a[31:29]};
            5'd30: y = { {30{sign}}, a[31:30]};
            5'd31: y = { {31{sign}}, a[31] };
            default: y = 32'b0;
        endcase
    end
endmodule

